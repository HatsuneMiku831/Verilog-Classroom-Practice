module decoder3_8( y,d );

    output [7:0] y;
    input [2:0] d;

    assign y[0] = ((~d[2]) & (~d[1]) & (~d[0])),
            y[1] = ((~d[2]) & (~d[1]) & (d[0])),
            y[2] = ((~d[2]) & (d[1]) & (~d[0])),
            y[3] = ((~d[2]) & (d[1]) & (d[0])),
            y[4] = ((d[2]) & (~d[1]) & (~d[0])),
            y[5] = ((d[2]) & (~d[1]) & (d[0])),
            y[6] = ((d[2]) & (d[1]) & (~d[0])),
            y[7] = ((d[2]) & (d[1]) & (d[0]));

endmodule